
package Sim6502_Package is

    type MemoryTransferType is (IDLE, READ, WRITE);

end package;
